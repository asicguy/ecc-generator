`timescale "1 ns / 10 ps"
