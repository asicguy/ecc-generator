////////////////////////////////////////////////////////////////
//
//  File name    : checker.sv
//  Creator      : Wang, Jun (phdbreak[at]gmail.com)
//
//  Results checker
// 
////////////////////////////////////////////////////////////////

`include "timescale.sv"
`include "define.sv"

program checker ();

// TODO

endprogram : checker
